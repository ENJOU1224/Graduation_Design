module HalfAdder (
	input		a,
	input		b,
	output	s	
);
	xor(s,a,b);
endmodule
